`timescale 1 ns / 10 ps

module convLayerMulti_TB();
parameter DATA_WIDTH = 16;
parameter D = 1; //Depth of image and filter
parameter H = 4; //Height of image
parameter W = 4; //Width of image
parameter F = 2; //Size of filter
parameter K = 1; //Number of filters applied
reg reset, clk;
reg [D*H*W*DATA_WIDTH-1:0] image;
reg [K*D*F*F*DATA_WIDTH-1:0] filters;
wire [0:K*(H-F+1)*(W-F+1)*DATA_WIDTH-1] outputConv;

localparam PERIOD = 100;

integer i;

always
	#(PERIOD/2) clk = ~clk;
	
	
initial begin 
	#0
	clk = 1'b0;
	reset = 1;
	//We test with a 1*32*32 image and 6 5*5 filters, all the values are 4
	//Expected output 4704 (6*28*28) values equal to 400 (16*25)
	image = 256'h3C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C00;
 	filters[0*F*F*DATA_WIDTH+:F*F*DATA_WIDTH] = 64'h3C003C003C003C00;
  	//filters[1*5*5*32+:5*5*32] = 800'h40800000408000004080000040800000408000004080000040800000408000004080000040800000408000004080000040800000408000004080000040800000408000004080000040800000408000004080000040800000408000004080000040800000;
  	//filters[2*5*5*32+:5*5*32] = 800'h40000000400000004000000040000000400000004000000040000000400000004000000040000000400000004000000040000000400000004000000040000000400000004000000040000000400000004000000040000000400000004000000040000000;	
  	//filters[3*5*5*32+:5*5*32] = 800'h40000000400000004000000040000000400000004000000040000000400000004000000040000000400000004000000040000000400000004000000040000000400000004000000040000000400000004000000040000000400000004000000040000000;	
  	//filters[4*5*5*32+:5*5*32] = 800'h40000000400000004000000040000000400000004000000040000000400000004000000040000000400000004000000040000000400000004000000040000000400000004000000040000000400000004000000040000000400000004000000040000000;	
  	//filters[5*5*5*32+:5*5*32] = 800'h40800000408000004080000040800000408000004080000040800000408000004080000040800000408000004080000040800000408000004080000040800000408000004080000040800000408000004080000040800000408000004080000040800000;

	#PERIOD
	reset = 0;

	
	#(((H-F+2)*(H-F)+1)*PERIOD)
	for (i = K*(H-F+1)*(H-F+1)-1; i >=0; i = i - 1) begin
		$displayh(outputConv[i*DATA_WIDTH+:DATA_WIDTH]);
	end
	$stop;
end

convLayerMulti #(
    .DATA_WIDTH ( DATA_WIDTH ),
    .D ( D ),
    .H ( H ),
    .W ( W ),
	.F ( F ),
    .K ( K )
)UUT(
	.clk(clk),
	.reset(reset),
	.image(image),
	.filters(filters),
	.outputConv(outputConv)
);

endmodule

