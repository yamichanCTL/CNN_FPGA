`timescale 100 ns / 10 ps

module convCal_TB #(
	parameter DATA_WIDTH = 16,
	parameter INPUT_CHANNEL = 2,
	parameter IMAGE_LENGTH = 4,
	parameter IMAGE_WIDTH = 4,

	parameter WEIGHT_LENGTH = 3,
	parameter WEIGHT_WIDTH = 3,
	parameter OUTPUT_CHANNEL = 2,

	parameter RESULT_LENGTH = 2,
	parameter RESULT_WIDTH = 2
)
();

reg clk, reset,conv_en;
reg [0:OUTPUT_CHANNEL*RESULT_LENGTH*RESULT_WIDTH*INPUT_CHANNEL*IMAGE_LENGTH*IMAGE_WIDTH*DATA_WIDTH-1] image;
reg [0:OUTPUT_CHANNEL*RESULT_LENGTH*RESULT_WIDTH*INPUT_CHANNEL*WEIGHT_LENGTH*WEIGHT_WIDTH*DATA_WIDTH-1] weight;

wire [0:OUTPUT_CHANNEL*RESULT_LENGTH*RESULT_WIDTH*DATA_WIDTH-1] result;
wire cc_valid;

localparam PERIOD = 2;

always
	#(PERIOD/2) clk = ~clk;

initial begin
	#0
	clk = 1'b0;reset = 1;conv_en = 0;
	// We test with an image part and a filter whose values are all 4 
	image =  4096'h3C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C00_3C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C00_3C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C00_3C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C00_3C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C00_3C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C00_3C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C00_3C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C00;
	weight=  2304'h3C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C00_3C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C00_3C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C00_3C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C00_3C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C00_3C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C00_3C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C00_3C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C003C00;
	
	#PERIOD reset = 0;conv_en = 1;

    #40 
	image =  4096'h40004000400040004000400040004000400040004000400040004000400040004000400040004000400040004000400040004000400040004000400040004000_40004000400040004000400040004000400040004000400040004000400040004000400040004000400040004000400040004000400040004000400040004000_40004000400040004000400040004000400040004000400040004000400040004000400040004000400040004000400040004000400040004000400040004000_40004000400040004000400040004000400040004000400040004000400040004000400040004000400040004000400040004000400040004000400040004000_40004000400040004000400040004000400040004000400040004000400040004000400040004000400040004000400040004000400040004000400040004000_40004000400040004000400040004000400040004000400040004000400040004000400040004000400040004000400040004000400040004000400040004000_40004000400040004000400040004000400040004000400040004000400040004000400040004000400040004000400040004000400040004000400040004000_40004000400040004000400040004000400040004000400040004000400040004000400040004000400040004000400040004000400040004000400040004000;
	//weight = 2304'h3C003C003C00_3C003C003C00_3C003C003C00_3C003C003C00_3C003C003C00_3C003C003C00;
	
end

convCal 
#(
	.DATA_WIDTH(DATA_WIDTH),
	.INPUT_CHANNEL(INPUT_CHANNEL),
	.IMAGE_LENGTH(IMAGE_LENGTH),
	.IMAGE_WIDTH(IMAGE_WIDTH),
    .WEIGHT_LENGTH(WEIGHT_LENGTH),
    .WEIGHT_WIDTH(WEIGHT_WIDTH),
    .OUTPUT_CHANNEL(OUTPUT_CHANNEL),
    .RESULT_LENGTH(RESULT_LENGTH),
    .RESULT_WIDTH(RESULT_WIDTH)
)
UUT
(
	.clk(clk),
	.reset(reset),
	.image(image),
	.conv_en(conv_en),
	.weight(weight),
	.result(result),
	.cc_valid(cc_valid)
);

endmodule
